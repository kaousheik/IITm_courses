module test_four_bit_adder;
reg [3:0] a,b;
reg s;

wire [4:0] sum2;
wire cout;

t3 DUT(a,b,s,sum2,cout);

initial
begin
$dumpfile("testfive.vcd");
$dumpvars(0,test_four_bit_adder);
$monitor("At time = %t, a  =  %b , b  =  %b  ,  s = %b , Output= %b",$time,a,b,s,sum2);
#10 a = 4'b0000; b = 4'b0000; s = 1'b0;
#10 a = 4'b0000; b = 4'b0001; s = 1'b0;
#10 a = 4'b0000; b = 4'b0010; s = 1'b0;
#10 a = 4'b0000; b = 4'b0011; s = 1'b0;
#10 a = 4'b0000; b = 4'b0100; s = 1'b0;
#10 a = 4'b0000; b = 4'b0101; s = 1'b0;
#10 a = 4'b0000; b = 4'b0110; s = 1'b0;
#10 a = 4'b0000; b = 4'b0111; s = 1'b0;
#10 a = 4'b0000; b = 4'b1000; s = 1'b0;
#10 a = 4'b0000; b = 4'b1001; s = 1'b0;
#10 a = 4'b0000; b = 4'b1010; s = 1'b0;
#10 a = 4'b0000; b = 4'b1011; s = 1'b0;
#10 a = 4'b0000; b = 4'b1100; s = 1'b0;
#10 a = 4'b0000; b = 4'b1101; s = 1'b0;
#10 a = 4'b0000; b = 4'b1110; s = 1'b0;
#10 a = 4'b0000; b = 4'b1111; s = 1'b0;
#10 a = 4'b0001; b = 4'b0000; s = 1'b0;
#10 a = 4'b0001; b = 4'b0001; s = 1'b0;
#10 a = 4'b0001; b = 4'b0010; s = 1'b0;
#10 a = 4'b0001; b = 4'b0011; s = 1'b0;
#10 a = 4'b0001; b = 4'b0100; s = 1'b0;
#10 a = 4'b0001; b = 4'b0101; s = 1'b0;
#10 a = 4'b0001; b = 4'b0110; s = 1'b0;
#10 a = 4'b0001; b = 4'b0111; s = 1'b0;
#10 a = 4'b0001; b = 4'b1000; s = 1'b0;
#10 a = 4'b0001; b = 4'b1001; s = 1'b0;
#10 a = 4'b0001; b = 4'b1010; s = 1'b0;
#10 a = 4'b0001; b = 4'b1011; s = 1'b0;
#10 a = 4'b0001; b = 4'b1100; s = 1'b0;
#10 a = 4'b0001; b = 4'b1101; s = 1'b0;
#10 a = 4'b0001; b = 4'b1110; s = 1'b0;
#10 a = 4'b0001; b = 4'b1111; s = 1'b0;
#10 a = 4'b0010; b = 4'b0000; s = 1'b0;
#10 a = 4'b0010; b = 4'b0001; s = 1'b0;
#10 a = 4'b0010; b = 4'b0010; s = 1'b0;
#10 a = 4'b0010; b = 4'b0011; s = 1'b0;
#10 a = 4'b0010; b = 4'b0100; s = 1'b0;
#10 a = 4'b0010; b = 4'b0101; s = 1'b0;
#10 a = 4'b0010; b = 4'b0110; s = 1'b0;
#10 a = 4'b0010; b = 4'b0111; s = 1'b0;
#10 a = 4'b0010; b = 4'b1000; s = 1'b0;
#10 a = 4'b0010; b = 4'b1001; s = 1'b0;
#10 a = 4'b0010; b = 4'b1010; s = 1'b0;
#10 a = 4'b0010; b = 4'b1011; s = 1'b0;
#10 a = 4'b0010; b = 4'b1100; s = 1'b0;
#10 a = 4'b0010; b = 4'b1101; s = 1'b0;
#10 a = 4'b0010; b = 4'b1110; s = 1'b0;
#10 a = 4'b0010; b = 4'b1111; s = 1'b0;
#10 a = 4'b0011; b = 4'b0000; s = 1'b0;
#10 a = 4'b0011; b = 4'b0001; s = 1'b0;
#10 a = 4'b0011; b = 4'b0010; s = 1'b0;
#10 a = 4'b0011; b = 4'b0011; s = 1'b0;
#10 a = 4'b0011; b = 4'b0100; s = 1'b0;
#10 a = 4'b0011; b = 4'b0101; s = 1'b0;
#10 a = 4'b0011; b = 4'b0110; s = 1'b0;
#10 a = 4'b0011; b = 4'b0111; s = 1'b0;
#10 a = 4'b0011; b = 4'b1000; s = 1'b0;
#10 a = 4'b0011; b = 4'b1001; s = 1'b0;
#10 a = 4'b0011; b = 4'b1010; s = 1'b0;
#10 a = 4'b0011; b = 4'b1011; s = 1'b0;
#10 a = 4'b0011; b = 4'b1100; s = 1'b0;
#10 a = 4'b0011; b = 4'b1101; s = 1'b0;
#10 a = 4'b0011; b = 4'b1110; s = 1'b0;
#10 a = 4'b0011; b = 4'b1111; s = 1'b0;
#10 a = 4'b0100; b = 4'b0000; s = 1'b0;
#10 a = 4'b0100; b = 4'b0001; s = 1'b0;
#10 a = 4'b0100; b = 4'b0010; s = 1'b0;
#10 a = 4'b0100; b = 4'b0011; s = 1'b0;
#10 a = 4'b0100; b = 4'b0100; s = 1'b0;
#10 a = 4'b0100; b = 4'b0101; s = 1'b0;
#10 a = 4'b0100; b = 4'b0110; s = 1'b0;
#10 a = 4'b0100; b = 4'b0111; s = 1'b0;
#10 a = 4'b0100; b = 4'b1000; s = 1'b0;
#10 a = 4'b0100; b = 4'b1001; s = 1'b0;
#10 a = 4'b0100; b = 4'b1010; s = 1'b0;
#10 a = 4'b0100; b = 4'b1011; s = 1'b0;
#10 a = 4'b0100; b = 4'b1100; s = 1'b0;
#10 a = 4'b0100; b = 4'b1101; s = 1'b0;
#10 a = 4'b0100; b = 4'b1110; s = 1'b0;
#10 a = 4'b0100; b = 4'b1111; s = 1'b0;
#10 a = 4'b0101; b = 4'b0000; s = 1'b0;
#10 a = 4'b0101; b = 4'b0001; s = 1'b0;
#10 a = 4'b0101; b = 4'b0010; s = 1'b0;
#10 a = 4'b0101; b = 4'b0011; s = 1'b0;
#10 a = 4'b0101; b = 4'b0100; s = 1'b0;
#10 a = 4'b0101; b = 4'b0101; s = 1'b0;
#10 a = 4'b0101; b = 4'b0110; s = 1'b0;
#10 a = 4'b0101; b = 4'b0111; s = 1'b0;
#10 a = 4'b0101; b = 4'b1000; s = 1'b0;
#10 a = 4'b0101; b = 4'b1001; s = 1'b0;
#10 a = 4'b0101; b = 4'b1010; s = 1'b0;
#10 a = 4'b0101; b = 4'b1011; s = 1'b0;
#10 a = 4'b0101; b = 4'b1100; s = 1'b0;
#10 a = 4'b0101; b = 4'b1101; s = 1'b0;
#10 a = 4'b0101; b = 4'b1110; s = 1'b0;
#10 a = 4'b0101; b = 4'b1111; s = 1'b0;
#10 a = 4'b0110; b = 4'b0000; s = 1'b0;
#10 a = 4'b0110; b = 4'b0001; s = 1'b0;
#10 a = 4'b0110; b = 4'b0010; s = 1'b0;
#10 a = 4'b0110; b = 4'b0011; s = 1'b0;
#10 a = 4'b0110; b = 4'b0100; s = 1'b0;
#10 a = 4'b0110; b = 4'b0101; s = 1'b0;
#10 a = 4'b0110; b = 4'b0110; s = 1'b0;
#10 a = 4'b0110; b = 4'b0111; s = 1'b0;
#10 a = 4'b0110; b = 4'b1000; s = 1'b0;
#10 a = 4'b0110; b = 4'b1001; s = 1'b0;
#10 a = 4'b0110; b = 4'b1010; s = 1'b0;
#10 a = 4'b0110; b = 4'b1011; s = 1'b0;
#10 a = 4'b0110; b = 4'b1100; s = 1'b0;
#10 a = 4'b0110; b = 4'b1101; s = 1'b0;
#10 a = 4'b0110; b = 4'b1110; s = 1'b0;
#10 a = 4'b0110; b = 4'b1111; s = 1'b0;
#10 a = 4'b0111; b = 4'b0000; s = 1'b0;
#10 a = 4'b0111; b = 4'b0001; s = 1'b0;
#10 a = 4'b0111; b = 4'b0010; s = 1'b0;
#10 a = 4'b0111; b = 4'b0011; s = 1'b0;
#10 a = 4'b0111; b = 4'b0100; s = 1'b0;
#10 a = 4'b0111; b = 4'b0101; s = 1'b0;
#10 a = 4'b0111; b = 4'b0110; s = 1'b0;
#10 a = 4'b0111; b = 4'b0111; s = 1'b0;
#10 a = 4'b0111; b = 4'b1000; s = 1'b0;
#10 a = 4'b0111; b = 4'b1001; s = 1'b0;
#10 a = 4'b0111; b = 4'b1010; s = 1'b0;
#10 a = 4'b0111; b = 4'b1011; s = 1'b0;
#10 a = 4'b0111; b = 4'b1100; s = 1'b0;
#10 a = 4'b0111; b = 4'b1101; s = 1'b0;
#10 a = 4'b0111; b = 4'b1110; s = 1'b0;
#10 a = 4'b0111; b = 4'b1111; s = 1'b0;
#10 a = 4'b1000; b = 4'b0000; s = 1'b0;
#10 a = 4'b1000; b = 4'b0001; s = 1'b0;
#10 a = 4'b1000; b = 4'b0010; s = 1'b0;
#10 a = 4'b1000; b = 4'b0011; s = 1'b0;
#10 a = 4'b1000; b = 4'b0100; s = 1'b0;
#10 a = 4'b1000; b = 4'b0101; s = 1'b0;
#10 a = 4'b1000; b = 4'b0110; s = 1'b0;
#10 a = 4'b1000; b = 4'b0111; s = 1'b0;
#10 a = 4'b1000; b = 4'b1000; s = 1'b0;
#10 a = 4'b1000; b = 4'b1001; s = 1'b0;
#10 a = 4'b1000; b = 4'b1010; s = 1'b0;
#10 a = 4'b1000; b = 4'b1011; s = 1'b0;
#10 a = 4'b1000; b = 4'b1100; s = 1'b0;
#10 a = 4'b1000; b = 4'b1101; s = 1'b0;
#10 a = 4'b1000; b = 4'b1110; s = 1'b0;
#10 a = 4'b1000; b = 4'b1111; s = 1'b0;
#10 a = 4'b1001; b = 4'b0000; s = 1'b0;
#10 a = 4'b1001; b = 4'b0001; s = 1'b0;
#10 a = 4'b1001; b = 4'b0010; s = 1'b0;
#10 a = 4'b1001; b = 4'b0011; s = 1'b0;
#10 a = 4'b1001; b = 4'b0100; s = 1'b0;
#10 a = 4'b1001; b = 4'b0101; s = 1'b0;
#10 a = 4'b1001; b = 4'b0110; s = 1'b0;
#10 a = 4'b1001; b = 4'b0111; s = 1'b0;
#10 a = 4'b1001; b = 4'b1000; s = 1'b0;
#10 a = 4'b1001; b = 4'b1001; s = 1'b0;
#10 a = 4'b1001; b = 4'b1010; s = 1'b0;
#10 a = 4'b1001; b = 4'b1011; s = 1'b0;
#10 a = 4'b1001; b = 4'b1100; s = 1'b0;
#10 a = 4'b1001; b = 4'b1101; s = 1'b0;
#10 a = 4'b1001; b = 4'b1110; s = 1'b0;
#10 a = 4'b1001; b = 4'b1111; s = 1'b0;
#10 a = 4'b1010; b = 4'b0000; s = 1'b0;
#10 a = 4'b1010; b = 4'b0001; s = 1'b0;
#10 a = 4'b1010; b = 4'b0010; s = 1'b0;
#10 a = 4'b1010; b = 4'b0011; s = 1'b0;
#10 a = 4'b1010; b = 4'b0100; s = 1'b0;
#10 a = 4'b1010; b = 4'b0101; s = 1'b0;
#10 a = 4'b1010; b = 4'b0110; s = 1'b0;
#10 a = 4'b1010; b = 4'b0111; s = 1'b0;
#10 a = 4'b1010; b = 4'b1000; s = 1'b0;
#10 a = 4'b1010; b = 4'b1001; s = 1'b0;
#10 a = 4'b1010; b = 4'b1010; s = 1'b0;
#10 a = 4'b1010; b = 4'b1011; s = 1'b0;
#10 a = 4'b1010; b = 4'b1100; s = 1'b0;
#10 a = 4'b1010; b = 4'b1101; s = 1'b0;
#10 a = 4'b1010; b = 4'b1110; s = 1'b0;
#10 a = 4'b1010; b = 4'b1111; s = 1'b0;
#10 a = 4'b1011; b = 4'b0000; s = 1'b0;
#10 a = 4'b1011; b = 4'b0001; s = 1'b0;
#10 a = 4'b1011; b = 4'b0010; s = 1'b0;
#10 a = 4'b1011; b = 4'b0011; s = 1'b0;
#10 a = 4'b1011; b = 4'b0100; s = 1'b0;
#10 a = 4'b1011; b = 4'b0101; s = 1'b0;
#10 a = 4'b1011; b = 4'b0110; s = 1'b0;
#10 a = 4'b1011; b = 4'b0111; s = 1'b0;
#10 a = 4'b1011; b = 4'b1000; s = 1'b0;
#10 a = 4'b1011; b = 4'b1001; s = 1'b0;
#10 a = 4'b1011; b = 4'b1010; s = 1'b0;
#10 a = 4'b1011; b = 4'b1011; s = 1'b0;
#10 a = 4'b1011; b = 4'b1100; s = 1'b0;
#10 a = 4'b1011; b = 4'b1101; s = 1'b0;
#10 a = 4'b1011; b = 4'b1110; s = 1'b0;
#10 a = 4'b1011; b = 4'b1111; s = 1'b0;
#10 a = 4'b1100; b = 4'b0000; s = 1'b0;
#10 a = 4'b1100; b = 4'b0001; s = 1'b0;
#10 a = 4'b1100; b = 4'b0010; s = 1'b0;
#10 a = 4'b1100; b = 4'b0011; s = 1'b0;
#10 a = 4'b1100; b = 4'b0100; s = 1'b0;
#10 a = 4'b1100; b = 4'b0101; s = 1'b0;
#10 a = 4'b1100; b = 4'b0110; s = 1'b0;
#10 a = 4'b1100; b = 4'b0111; s = 1'b0;
#10 a = 4'b1100; b = 4'b1000; s = 1'b0;
#10 a = 4'b1100; b = 4'b1001; s = 1'b0;
#10 a = 4'b1100; b = 4'b1010; s = 1'b0;
#10 a = 4'b1100; b = 4'b1011; s = 1'b0;
#10 a = 4'b1100; b = 4'b1100; s = 1'b0;
#10 a = 4'b1100; b = 4'b1101; s = 1'b0;
#10 a = 4'b1100; b = 4'b1110; s = 1'b0;
#10 a = 4'b1100; b = 4'b1111; s = 1'b0;
#10 a = 4'b1101; b = 4'b0000; s = 1'b0;
#10 a = 4'b1101; b = 4'b0001; s = 1'b0;
#10 a = 4'b1101; b = 4'b0010; s = 1'b0;
#10 a = 4'b1101; b = 4'b0011; s = 1'b0;
#10 a = 4'b1101; b = 4'b0100; s = 1'b0;
#10 a = 4'b1101; b = 4'b0101; s = 1'b0;
#10 a = 4'b1101; b = 4'b0110; s = 1'b0;
#10 a = 4'b1101; b = 4'b0111; s = 1'b0;
#10 a = 4'b1101; b = 4'b1000; s = 1'b0;
#10 a = 4'b1101; b = 4'b1001; s = 1'b0;
#10 a = 4'b1101; b = 4'b1010; s = 1'b0;
#10 a = 4'b1101; b = 4'b1011; s = 1'b0;
#10 a = 4'b1101; b = 4'b1100; s = 1'b0;
#10 a = 4'b1101; b = 4'b1101; s = 1'b0;
#10 a = 4'b1101; b = 4'b1110; s = 1'b0;
#10 a = 4'b1101; b = 4'b1111; s = 1'b0;
#10 a = 4'b1110; b = 4'b0000; s = 1'b0;
#10 a = 4'b1110; b = 4'b0001; s = 1'b0;
#10 a = 4'b1110; b = 4'b0010; s = 1'b0;
#10 a = 4'b1110; b = 4'b0011; s = 1'b0;
#10 a = 4'b1110; b = 4'b0100; s = 1'b0;
#10 a = 4'b1110; b = 4'b0101; s = 1'b0;
#10 a = 4'b1110; b = 4'b0110; s = 1'b0;
#10 a = 4'b1110; b = 4'b0111; s = 1'b0;
#10 a = 4'b1110; b = 4'b1000; s = 1'b0;
#10 a = 4'b1110; b = 4'b1001; s = 1'b0;
#10 a = 4'b1110; b = 4'b1010; s = 1'b0;
#10 a = 4'b1110; b = 4'b1011; s = 1'b0;
#10 a = 4'b1110; b = 4'b1100; s = 1'b0;
#10 a = 4'b1110; b = 4'b1101; s = 1'b0;
#10 a = 4'b1110; b = 4'b1110; s = 1'b0;
#10 a = 4'b1110; b = 4'b1111; s = 1'b0;
#10 a = 4'b1111; b = 4'b0000; s = 1'b0;
#10 a = 4'b1111; b = 4'b0001; s = 1'b0;
#10 a = 4'b1111; b = 4'b0010; s = 1'b0;
#10 a = 4'b1111; b = 4'b0011; s = 1'b0;
#10 a = 4'b1111; b = 4'b0100; s = 1'b0;
#10 a = 4'b1111; b = 4'b0101; s = 1'b0;
#10 a = 4'b1111; b = 4'b0110; s = 1'b0;
#10 a = 4'b1111; b = 4'b0111; s = 1'b0;
#10 a = 4'b1111; b = 4'b1000; s = 1'b0;
#10 a = 4'b1111; b = 4'b1001; s = 1'b0;
#10 a = 4'b1111; b = 4'b1010; s = 1'b0;
#10 a = 4'b1111; b = 4'b1011; s = 1'b0;
#10 a = 4'b1111; b = 4'b1100; s = 1'b0;
#10 a = 4'b1111; b = 4'b1101; s = 1'b0;
#10 a = 4'b1111; b = 4'b1110; s = 1'b0;
#10 a = 4'b1111; b = 4'b1111; s = 1'b0;
#10 a = 4'b0000; b = 4'b0000; s = 1'b1;
#10 a = 4'b0000; b = 4'b0001; s = 1'b1;
#10 a = 4'b0000; b = 4'b0010; s = 1'b1;
#10 a = 4'b0000; b = 4'b0011; s = 1'b1;
#10 a = 4'b0000; b = 4'b0100; s = 1'b1;
#10 a = 4'b0000; b = 4'b0101; s = 1'b1;
#10 a = 4'b0000; b = 4'b0110; s = 1'b1;
#10 a = 4'b0000; b = 4'b0111; s = 1'b1;
#10 a = 4'b0000; b = 4'b1000; s = 1'b1;
#10 a = 4'b0000; b = 4'b1001; s = 1'b1;
#10 a = 4'b0000; b = 4'b1010; s = 1'b1;
#10 a = 4'b0000; b = 4'b1011; s = 1'b1;
#10 a = 4'b0000; b = 4'b1100; s = 1'b1;
#10 a = 4'b0000; b = 4'b1101; s = 1'b1;
#10 a = 4'b0000; b = 4'b1110; s = 1'b1;
#10 a = 4'b0000; b = 4'b1111; s = 1'b1;
#10 a = 4'b0001; b = 4'b0000; s = 1'b1;
#10 a = 4'b0001; b = 4'b0001; s = 1'b1;
#10 a = 4'b0001; b = 4'b0010; s = 1'b1;
#10 a = 4'b0001; b = 4'b0011; s = 1'b1;
#10 a = 4'b0001; b = 4'b0100; s = 1'b1;
#10 a = 4'b0001; b = 4'b0101; s = 1'b1;
#10 a = 4'b0001; b = 4'b0110; s = 1'b1;
#10 a = 4'b0001; b = 4'b0111; s = 1'b1;
#10 a = 4'b0001; b = 4'b1000; s = 1'b1;
#10 a = 4'b0001; b = 4'b1001; s = 1'b1;
#10 a = 4'b0001; b = 4'b1010; s = 1'b1;
#10 a = 4'b0001; b = 4'b1011; s = 1'b1;
#10 a = 4'b0001; b = 4'b1100; s = 1'b1;
#10 a = 4'b0001; b = 4'b1101; s = 1'b1;
#10 a = 4'b0001; b = 4'b1110; s = 1'b1;
#10 a = 4'b0001; b = 4'b1111; s = 1'b1;
#10 a = 4'b0010; b = 4'b0000; s = 1'b1;
#10 a = 4'b0010; b = 4'b0001; s = 1'b1;
#10 a = 4'b0010; b = 4'b0010; s = 1'b1;
#10 a = 4'b0010; b = 4'b0011; s = 1'b1;
#10 a = 4'b0010; b = 4'b0100; s = 1'b1;
#10 a = 4'b0010; b = 4'b0101; s = 1'b1;
#10 a = 4'b0010; b = 4'b0110; s = 1'b1;
#10 a = 4'b0010; b = 4'b0111; s = 1'b1;
#10 a = 4'b0010; b = 4'b1000; s = 1'b1;
#10 a = 4'b0010; b = 4'b1001; s = 1'b1;
#10 a = 4'b0010; b = 4'b1010; s = 1'b1;
#10 a = 4'b0010; b = 4'b1011; s = 1'b1;
#10 a = 4'b0010; b = 4'b1100; s = 1'b1;
#10 a = 4'b0010; b = 4'b1101; s = 1'b1;
#10 a = 4'b0010; b = 4'b1110; s = 1'b1;
#10 a = 4'b0010; b = 4'b1111; s = 1'b1;
#10 a = 4'b0011; b = 4'b0000; s = 1'b1;
#10 a = 4'b0011; b = 4'b0001; s = 1'b1;
#10 a = 4'b0011; b = 4'b0010; s = 1'b1;
#10 a = 4'b0011; b = 4'b0011; s = 1'b1;
#10 a = 4'b0011; b = 4'b0100; s = 1'b1;
#10 a = 4'b0011; b = 4'b0101; s = 1'b1;
#10 a = 4'b0011; b = 4'b0110; s = 1'b1;
#10 a = 4'b0011; b = 4'b0111; s = 1'b1;
#10 a = 4'b0011; b = 4'b1000; s = 1'b1;
#10 a = 4'b0011; b = 4'b1001; s = 1'b1;
#10 a = 4'b0011; b = 4'b1010; s = 1'b1;
#10 a = 4'b0011; b = 4'b1011; s = 1'b1;
#10 a = 4'b0011; b = 4'b1100; s = 1'b1;
#10 a = 4'b0011; b = 4'b1101; s = 1'b1;
#10 a = 4'b0011; b = 4'b1110; s = 1'b1;
#10 a = 4'b0011; b = 4'b1111; s = 1'b1;
#10 a = 4'b0100; b = 4'b0000; s = 1'b1;
#10 a = 4'b0100; b = 4'b0001; s = 1'b1;
#10 a = 4'b0100; b = 4'b0010; s = 1'b1;
#10 a = 4'b0100; b = 4'b0011; s = 1'b1;
#10 a = 4'b0100; b = 4'b0100; s = 1'b1;
#10 a = 4'b0100; b = 4'b0101; s = 1'b1;
#10 a = 4'b0100; b = 4'b0110; s = 1'b1;
#10 a = 4'b0100; b = 4'b0111; s = 1'b1;
#10 a = 4'b0100; b = 4'b1000; s = 1'b1;
#10 a = 4'b0100; b = 4'b1001; s = 1'b1;
#10 a = 4'b0100; b = 4'b1010; s = 1'b1;
#10 a = 4'b0100; b = 4'b1011; s = 1'b1;
#10 a = 4'b0100; b = 4'b1100; s = 1'b1;
#10 a = 4'b0100; b = 4'b1101; s = 1'b1;
#10 a = 4'b0100; b = 4'b1110; s = 1'b1;
#10 a = 4'b0100; b = 4'b1111; s = 1'b1;
#10 a = 4'b0101; b = 4'b0000; s = 1'b1;
#10 a = 4'b0101; b = 4'b0001; s = 1'b1;
#10 a = 4'b0101; b = 4'b0010; s = 1'b1;
#10 a = 4'b0101; b = 4'b0011; s = 1'b1;
#10 a = 4'b0101; b = 4'b0100; s = 1'b1;
#10 a = 4'b0101; b = 4'b0101; s = 1'b1;
#10 a = 4'b0101; b = 4'b0110; s = 1'b1;
#10 a = 4'b0101; b = 4'b0111; s = 1'b1;
#10 a = 4'b0101; b = 4'b1000; s = 1'b1;
#10 a = 4'b0101; b = 4'b1001; s = 1'b1;
#10 a = 4'b0101; b = 4'b1010; s = 1'b1;
#10 a = 4'b0101; b = 4'b1011; s = 1'b1;
#10 a = 4'b0101; b = 4'b1100; s = 1'b1;
#10 a = 4'b0101; b = 4'b1101; s = 1'b1;
#10 a = 4'b0101; b = 4'b1110; s = 1'b1;
#10 a = 4'b0101; b = 4'b1111; s = 1'b1;
#10 a = 4'b0110; b = 4'b0000; s = 1'b1;
#10 a = 4'b0110; b = 4'b0001; s = 1'b1;
#10 a = 4'b0110; b = 4'b0010; s = 1'b1;
#10 a = 4'b0110; b = 4'b0011; s = 1'b1;
#10 a = 4'b0110; b = 4'b0100; s = 1'b1;
#10 a = 4'b0110; b = 4'b0101; s = 1'b1;
#10 a = 4'b0110; b = 4'b0110; s = 1'b1;
#10 a = 4'b0110; b = 4'b0111; s = 1'b1;
#10 a = 4'b0110; b = 4'b1000; s = 1'b1;
#10 a = 4'b0110; b = 4'b1001; s = 1'b1;
#10 a = 4'b0110; b = 4'b1010; s = 1'b1;
#10 a = 4'b0110; b = 4'b1011; s = 1'b1;
#10 a = 4'b0110; b = 4'b1100; s = 1'b1;
#10 a = 4'b0110; b = 4'b1101; s = 1'b1;
#10 a = 4'b0110; b = 4'b1110; s = 1'b1;
#10 a = 4'b0110; b = 4'b1111; s = 1'b1;
#10 a = 4'b0111; b = 4'b0000; s = 1'b1;
#10 a = 4'b0111; b = 4'b0001; s = 1'b1;
#10 a = 4'b0111; b = 4'b0010; s = 1'b1;
#10 a = 4'b0111; b = 4'b0011; s = 1'b1;
#10 a = 4'b0111; b = 4'b0100; s = 1'b1;
#10 a = 4'b0111; b = 4'b0101; s = 1'b1;
#10 a = 4'b0111; b = 4'b0110; s = 1'b1;
#10 a = 4'b0111; b = 4'b0111; s = 1'b1;
#10 a = 4'b0111; b = 4'b1000; s = 1'b1;
#10 a = 4'b0111; b = 4'b1001; s = 1'b1;
#10 a = 4'b0111; b = 4'b1010; s = 1'b1;
#10 a = 4'b0111; b = 4'b1011; s = 1'b1;
#10 a = 4'b0111; b = 4'b1100; s = 1'b1;
#10 a = 4'b0111; b = 4'b1101; s = 1'b1;
#10 a = 4'b0111; b = 4'b1110; s = 1'b1;
#10 a = 4'b0111; b = 4'b1111; s = 1'b1;
#10 a = 4'b1000; b = 4'b0000; s = 1'b1;
#10 a = 4'b1000; b = 4'b0001; s = 1'b1;
#10 a = 4'b1000; b = 4'b0010; s = 1'b1;
#10 a = 4'b1000; b = 4'b0011; s = 1'b1;
#10 a = 4'b1000; b = 4'b0100; s = 1'b1;
#10 a = 4'b1000; b = 4'b0101; s = 1'b1;
#10 a = 4'b1000; b = 4'b0110; s = 1'b1;
#10 a = 4'b1000; b = 4'b0111; s = 1'b1;
#10 a = 4'b1000; b = 4'b1000; s = 1'b1;
#10 a = 4'b1000; b = 4'b1001; s = 1'b1;
#10 a = 4'b1000; b = 4'b1010; s = 1'b1;
#10 a = 4'b1000; b = 4'b1011; s = 1'b1;
#10 a = 4'b1000; b = 4'b1100; s = 1'b1;
#10 a = 4'b1000; b = 4'b1101; s = 1'b1;
#10 a = 4'b1000; b = 4'b1110; s = 1'b1;
#10 a = 4'b1000; b = 4'b1111; s = 1'b1;
#10 a = 4'b1001; b = 4'b0000; s = 1'b1;
#10 a = 4'b1001; b = 4'b0001; s = 1'b1;
#10 a = 4'b1001; b = 4'b0010; s = 1'b1;
#10 a = 4'b1001; b = 4'b0011; s = 1'b1;
#10 a = 4'b1001; b = 4'b0100; s = 1'b1;
#10 a = 4'b1001; b = 4'b0101; s = 1'b1;
#10 a = 4'b1001; b = 4'b0110; s = 1'b1;
#10 a = 4'b1001; b = 4'b0111; s = 1'b1;
#10 a = 4'b1001; b = 4'b1000; s = 1'b1;
#10 a = 4'b1001; b = 4'b1001; s = 1'b1;
#10 a = 4'b1001; b = 4'b1010; s = 1'b1;
#10 a = 4'b1001; b = 4'b1011; s = 1'b1;
#10 a = 4'b1001; b = 4'b1100; s = 1'b1;
#10 a = 4'b1001; b = 4'b1101; s = 1'b1;
#10 a = 4'b1001; b = 4'b1110; s = 1'b1;
#10 a = 4'b1001; b = 4'b1111; s = 1'b1;
#10 a = 4'b1010; b = 4'b0000; s = 1'b1;
#10 a = 4'b1010; b = 4'b0001; s = 1'b1;
#10 a = 4'b1010; b = 4'b0010; s = 1'b1;
#10 a = 4'b1010; b = 4'b0011; s = 1'b1;
#10 a = 4'b1010; b = 4'b0100; s = 1'b1;
#10 a = 4'b1010; b = 4'b0101; s = 1'b1;
#10 a = 4'b1010; b = 4'b0110; s = 1'b1;
#10 a = 4'b1010; b = 4'b0111; s = 1'b1;
#10 a = 4'b1010; b = 4'b1000; s = 1'b1;
#10 a = 4'b1010; b = 4'b1001; s = 1'b1;
#10 a = 4'b1010; b = 4'b1010; s = 1'b1;
#10 a = 4'b1010; b = 4'b1011; s = 1'b1;
#10 a = 4'b1010; b = 4'b1100; s = 1'b1;
#10 a = 4'b1010; b = 4'b1101; s = 1'b1;
#10 a = 4'b1010; b = 4'b1110; s = 1'b1;
#10 a = 4'b1010; b = 4'b1111; s = 1'b1;
#10 a = 4'b1011; b = 4'b0000; s = 1'b1;
#10 a = 4'b1011; b = 4'b0001; s = 1'b1;
#10 a = 4'b1011; b = 4'b0010; s = 1'b1;
#10 a = 4'b1011; b = 4'b0011; s = 1'b1;
#10 a = 4'b1011; b = 4'b0100; s = 1'b1;
#10 a = 4'b1011; b = 4'b0101; s = 1'b1;
#10 a = 4'b1011; b = 4'b0110; s = 1'b1;
#10 a = 4'b1011; b = 4'b0111; s = 1'b1;
#10 a = 4'b1011; b = 4'b1000; s = 1'b1;
#10 a = 4'b1011; b = 4'b1001; s = 1'b1;
#10 a = 4'b1011; b = 4'b1010; s = 1'b1;
#10 a = 4'b1011; b = 4'b1011; s = 1'b1;
#10 a = 4'b1011; b = 4'b1100; s = 1'b1;
#10 a = 4'b1011; b = 4'b1101; s = 1'b1;
#10 a = 4'b1011; b = 4'b1110; s = 1'b1;
#10 a = 4'b1011; b = 4'b1111; s = 1'b1;
#10 a = 4'b1100; b = 4'b0000; s = 1'b1;
#10 a = 4'b1100; b = 4'b0001; s = 1'b1;
#10 a = 4'b1100; b = 4'b0010; s = 1'b1;
#10 a = 4'b1100; b = 4'b0011; s = 1'b1;
#10 a = 4'b1100; b = 4'b0100; s = 1'b1;
#10 a = 4'b1100; b = 4'b0101; s = 1'b1;
#10 a = 4'b1100; b = 4'b0110; s = 1'b1;
#10 a = 4'b1100; b = 4'b0111; s = 1'b1;
#10 a = 4'b1100; b = 4'b1000; s = 1'b1;
#10 a = 4'b1100; b = 4'b1001; s = 1'b1;
#10 a = 4'b1100; b = 4'b1010; s = 1'b1;
#10 a = 4'b1100; b = 4'b1011; s = 1'b1;
#10 a = 4'b1100; b = 4'b1100; s = 1'b1;
#10 a = 4'b1100; b = 4'b1101; s = 1'b1;
#10 a = 4'b1100; b = 4'b1110; s = 1'b1;
#10 a = 4'b1100; b = 4'b1111; s = 1'b1;
#10 a = 4'b1101; b = 4'b0000; s = 1'b1;
#10 a = 4'b1101; b = 4'b0001; s = 1'b1;
#10 a = 4'b1101; b = 4'b0010; s = 1'b1;
#10 a = 4'b1101; b = 4'b0011; s = 1'b1;
#10 a = 4'b1101; b = 4'b0100; s = 1'b1;
#10 a = 4'b1101; b = 4'b0101; s = 1'b1;
#10 a = 4'b1101; b = 4'b0110; s = 1'b1;
#10 a = 4'b1101; b = 4'b0111; s = 1'b1;
#10 a = 4'b1101; b = 4'b1000; s = 1'b1;
#10 a = 4'b1101; b = 4'b1001; s = 1'b1;
#10 a = 4'b1101; b = 4'b1010; s = 1'b1;
#10 a = 4'b1101; b = 4'b1011; s = 1'b1;
#10 a = 4'b1101; b = 4'b1100; s = 1'b1;
#10 a = 4'b1101; b = 4'b1101; s = 1'b1;
#10 a = 4'b1101; b = 4'b1110; s = 1'b1;
#10 a = 4'b1101; b = 4'b1111; s = 1'b1;
#10 a = 4'b1110; b = 4'b0000; s = 1'b1;
#10 a = 4'b1110; b = 4'b0001; s = 1'b1;
#10 a = 4'b1110; b = 4'b0010; s = 1'b1;
#10 a = 4'b1110; b = 4'b0011; s = 1'b1;
#10 a = 4'b1110; b = 4'b0100; s = 1'b1;
#10 a = 4'b1110; b = 4'b0101; s = 1'b1;
#10 a = 4'b1110; b = 4'b0110; s = 1'b1;
#10 a = 4'b1110; b = 4'b0111; s = 1'b1;
#10 a = 4'b1110; b = 4'b1000; s = 1'b1;
#10 a = 4'b1110; b = 4'b1001; s = 1'b1;
#10 a = 4'b1110; b = 4'b1010; s = 1'b1;
#10 a = 4'b1110; b = 4'b1011; s = 1'b1;
#10 a = 4'b1110; b = 4'b1100; s = 1'b1;
#10 a = 4'b1110; b = 4'b1101; s = 1'b1;
#10 a = 4'b1110; b = 4'b1110; s = 1'b1;
#10 a = 4'b1110; b = 4'b1111; s = 1'b1;
#10 a = 4'b1111; b = 4'b0000; s = 1'b1;
#10 a = 4'b1111; b = 4'b0001; s = 1'b1;
#10 a = 4'b1111; b = 4'b0010; s = 1'b1;
#10 a = 4'b1111; b = 4'b0011; s = 1'b1;
#10 a = 4'b1111; b = 4'b0100; s = 1'b1;
#10 a = 4'b1111; b = 4'b0101; s = 1'b1;
#10 a = 4'b1111; b = 4'b0110; s = 1'b1;
#10 a = 4'b1111; b = 4'b0111; s = 1'b1;
#10 a = 4'b1111; b = 4'b1000; s = 1'b1;
#10 a = 4'b1111; b = 4'b1001; s = 1'b1;
#10 a = 4'b1111; b = 4'b1010; s = 1'b1;
#10 a = 4'b1111; b = 4'b1011; s = 1'b1;
#10 a = 4'b1111; b = 4'b1100; s = 1'b1;
#10 a = 4'b1111; b = 4'b1101; s = 1'b1;
#10 a = 4'b1111; b = 4'b1110; s = 1'b1;
#10 a = 4'b1111; b = 4'b1111; s = 1'b1;

#10 $finish;
end
endmodule
